module Processador

endmodule
